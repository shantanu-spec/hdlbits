module top_module (
    input [31:0] a,
    input [31:0] b,
    output [31:0] sum
);//
    wire temp,temp2;
    add16 adder1(a[15:0],b[15:0],0,sum[15:0],temp);
    add16 adder2(a[31:16],b[31:16],temp,sum[31:16],temp2);
    
endmodule

module add1 ( input a, input b, input cin,   output sum, output cout );
 assign {cout, sum} = a + b + cin;
// Full adder module here

endmodule
